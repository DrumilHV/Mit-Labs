module q1(W,F);
    input [3:0]W;
    // input En;
    // output [15:0]Y;
    output F;
    wire [0:15]Y;
    dec4to16 dec(W,Y);
    assign F = Y[1] | Y[3] | Y[6] | Y[7] | Y[9] | Y[14] | Y[15];
endmodule

module dec4to16(W,Y);
    input [3:0]W;
    // input En;
    output [15:0]Y;
    reg [15:0]Y;
    always@(W)
    begin
        // if(En==0)
            // Y=16'b0000000000000000;
        // else
            case(W)
                0:Y=16'b1000000000000000;
                1:Y=16'b0100000000000000;
                2:Y=16'b0010000000000000;
                3:Y=16'b0001000000000000;
                4:Y=16'b0000100000000000;
                5:Y=16'b0000010000000000;
                6:Y=16'b0000001000000000;
                7:Y=16'b0000000100000000;
                8:Y=16'b0000000010000000;
                9:Y=16'b0000000001000000;
                10:Y=16'b000000000100000;
                11:Y=16'b000000000010000;
                12:Y=16'b000000000001000;
                13:Y=16'b000000000000100;
                14:Y=16'b000000000000010;
                15:Y=16'b000000000000001;
            endcase
    end
endmodule
